module Lab9(clk, rst, ALUout, instr, immSel, regRW, ALUsrc, ALUop, MRW, PCsrc, WB, ALU1, readRS1, readRS2, currentPC, nextPC, immOut, offsetPC, writeRD, dataOut);

	input clk, rst;
	
	// Test outputs
	output [31:0] ALUout, ALU1, readRS1, readRS2, currentPC, nextPC, immOut, offsetPC, writeRD, dataOut;
	output [31:0] instr;
	output [1:0] immSel;
	output [1:0] regRW;
	output ALUsrc;
	output [3:0] ALUop;
	output MRW;
	output PCsrc;
	output WB;
	
	// Datapath / Control Unit Interconnects
	wire [31:0] instr;
	wire [1:0] immSel;
	wire [1:0] regRW;
	wire ALUsrc;
	wire [1:0] status;
	wire [2:0] ALUop;
	wire MRW;
	wire PCsrc;
	wire WB;
	
	ControlUnit CU(clk, rst, instr, immSel, regRW, ALUsrc, status, ALUop, MRW, PCsrc, WB);
	
	Datapath DP(clk, rst, instr, immSel, regRW, ALUsrc, status, ALUop, MRW, PCsrc, WB, readRS1, ALU1, ALUout, readRS2, dataOut, currentPC, nextPC, immOut, offsetPC, writeRD);
	

endmodule
